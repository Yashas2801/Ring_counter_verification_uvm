package ring_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "ring_xtn.sv"

  `include "ring_seqs.sv"

  `include "ring_driver.sv"
  `include "ring_monitor.sv"
  `include "ring_sequencer.sv"
  `include "ring_agent.sv"

  `include "ring_coverage.sv"
  `include "ring_env.sv"

  `include "ring_test.sv"
endpackage
